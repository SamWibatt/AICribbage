.title KiCad schematic
P8 NC_01 CONN_01X01
P9 NC_02 CONN_01X01
P10 NC_03 CONN_01X01
P11 NC_04 CONN_01X01
P12 NC_05 CONN_01X01
P13 NC_06 CONN_01X01
P2 NC_07 NC_08 NC_09 +3V3 +5V GND GND NC_10 Power
P5 NC_11 NC_12 NC_13 GND /13_**_ /12_**_ /11_**_ /10_**_ /9_**_ /8_**_ PWM
P6 /7_**_ /6_**_ /5_**_ /4_**_ /3_**_ /2_**_ /1_Tx0_ /0_Rx0_ PWM
P4 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 Analog
P7 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 Communication
P1 GND GND NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 NC_51 NC_52 NC_53 NC_54 NC_55 NC_56 NC_57 NC_58 NC_59 NC_60 NC_61 +5V +5V Digital
U1 NC_62 NC_63 /A0 NC_64 NC_65 NC_66 /A1 /A2 /A3 /A4 /8_**_ /9_**_ /4_**_ /3_**_ /1_Tx0_ /0_Rx0_ NC_67 NC_68 NC_69 NC_70 NC_71 NC_72 /2_**_ /5_**_ /11_**_ /13_**_ /10_**_ /12_**_ /6_**_ /7_**_ NC_73 NC_74 NC_75 NC_76 NC_77 NC_78 NC_79 NC_80 NC_81 NC_82 NC_83 NC_84 NC_85 NC_86 NC_87 NC_88 /A5 NC_89 NC_90 ATSAMD21G18A-AU
U2 NC_91 NC_92 NC_93 L7805
P3 /A0 /A1 /A2 /A3 /A4 /A5 NC_94 NC_95 Analog
.end
